module m;
    // hello
    bit [4:0] b;
    int b;
    begin end
endmodule