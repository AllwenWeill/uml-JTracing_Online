module m;
    // hello
    bit [4:0] b;
    int b; //注意：此处有重命名错误
    begin end
endmodule