reg [0:1] port;
parameter a = 5;
module m;
____________________
module m(
    input port1 a;
    output port2 b;
)