int a = 0;
for (int i = 0; i <= 5; i++) begin
        a = a + 1;
end