module m;
    // hello
    string s = "hello world";
    begin end
endmodule