module m;
    // hello
    string s = "FOO";

    begin end
endmodule

